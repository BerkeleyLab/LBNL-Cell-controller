localparam QSFP1_VENDOR_NAME = 'h0;
localparam QSFP1_VENDOR_NAME_SIZE = 16;
localparam QSFP1_PART_NAME = 'h10;
localparam QSFP1_PART_NAME_SIZE = 16;
localparam QSFP1_REVISION_CODE = 'h20;
localparam QSFP1_REVISION_CODE_SIZE = 2;
localparam QSFP1_WAVELENGTH = 'h22;
localparam QSFP1_WAVELENGTH_SIZE = 2;
localparam QSFP1_SER_NUM = 'h24;
localparam QSFP1_SER_NUM_SIZE = 16;
localparam QSFP1_DATE_CODE = 'h34;
localparam QSFP1_DATE_CODE_SIZE = 8;
localparam QSFP2_VENDOR_NAME = 'h3c;
localparam QSFP2_VENDOR_NAME_SIZE = 16;
localparam QSFP2_PART_NAME = 'h4c;
localparam QSFP2_PART_NAME_SIZE = 16;
localparam QSFP2_REVISION_CODE = 'h5c;
localparam QSFP2_REVISION_CODE_SIZE = 2;
localparam QSFP2_WAVELENGTH = 'h5e;
localparam QSFP2_WAVELENGTH_SIZE = 2;
localparam QSFP2_SER_NUM = 'h60;
localparam QSFP2_SER_NUM_SIZE = 16;
localparam QSFP2_DATE_CODE = 'h70;
localparam QSFP2_DATE_CODE_SIZE = 8;
localparam U34_PORT_DATA = 'h80;
localparam U34_PORT_DATA_SIZE = 2;
localparam U39_PORT_DATA = 'h82;
localparam U39_PORT_DATA_SIZE = 2;
localparam QSFP1_MODULE_STATUS = 'h84;
localparam QSFP1_MODULE_STATUS_SIZE = 1;
localparam QSFP1_TEMPERATURE = 'h85;
localparam QSFP1_TEMPERATURE_SIZE = 2;
localparam QSFP1_VSUPPLY = 'h87;
localparam QSFP1_VSUPPLY_SIZE = 2;
localparam QSFP1_RXPOWER = 'h89;
localparam QSFP1_RXPOWER_SIZE = 8;
localparam QSFP1_IDENTIFIER = 'h91;
localparam QSFP1_IDENTIFIER_SIZE = 2;
localparam QSFP2_MODULE_STATUS = 'h93;
localparam QSFP2_MODULE_STATUS_SIZE = 1;
localparam QSFP2_TEMPERATURE = 'h94;
localparam QSFP2_TEMPERATURE_SIZE = 2;
localparam QSFP2_VSUPPLY = 'h96;
localparam QSFP2_VSUPPLY_SIZE = 2;
localparam QSFP2_RXPOWER = 'h98;
localparam QSFP2_RXPOWER_SIZE = 8;
localparam QSFP2_IDENTIFIER = 'ha0;
localparam QSFP2_IDENTIFIER_SIZE = 2;
