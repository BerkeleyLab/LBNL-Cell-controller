localparam QSFP1_VENDOR_NAME = 'h0;
localparam QSFP1_VENDOR_NAME_SIZE = 16;
localparam QSFP1_PART_NAME = 'h10;
localparam QSFP1_PART_NAME_SIZE = 16;
localparam QSFP1_REVISION_CODE = 'h20;
localparam QSFP1_REVISION_CODE_SIZE = 2;
localparam QSFP1_WAVELENGTH = 'h22;
localparam QSFP1_WAVELENGTH_SIZE = 2;
localparam QSFP1_SER_NUM = 'h24;
localparam QSFP1_SER_NUM_SIZE = 16;
localparam QSFP1_DATE_CODE = 'h34;
localparam QSFP1_DATE_CODE_SIZE = 8;
localparam QSFP2_VENDOR_NAME = 'h3c;
localparam QSFP2_VENDOR_NAME_SIZE = 16;
localparam QSFP2_PART_NAME = 'h4c;
localparam QSFP2_PART_NAME_SIZE = 16;
localparam QSFP2_REVISION_CODE = 'h5c;
localparam QSFP2_REVISION_CODE_SIZE = 2;
localparam QSFP2_WAVELENGTH = 'h5e;
localparam QSFP2_WAVELENGTH_SIZE = 2;
localparam QSFP2_SER_NUM = 'h60;
localparam QSFP2_SER_NUM_SIZE = 16;
localparam QSFP2_DATE_CODE = 'h70;
localparam QSFP2_DATE_CODE_SIZE = 8;
localparam U34_PORT0 = 'h78;
localparam U34_PORT0_SIZE = 1;
localparam U34_PORT1 = 'h79;
localparam U34_PORT1_SIZE = 1;
localparam QSFP1_MODULE_STATUS = 'h7a;
localparam QSFP1_MODULE_STATUS_SIZE = 1;
localparam QSFP1_TEMPERATURE = 'h7b;
localparam QSFP1_TEMPERATURE_SIZE = 2;
localparam QSFP1_VSUPPLY = 'h7d;
localparam QSFP1_VSUPPLY_SIZE = 2;
localparam QSFP1_RXPOWER = 'h7f;
localparam QSFP1_RXPOWER_SIZE = 8;
localparam QSFP1_IDENTIFIER = 'h87;
localparam QSFP1_IDENTIFIER_SIZE = 2;
localparam QSFP2_MODULE_STATUS = 'h89;
localparam QSFP2_MODULE_STATUS_SIZE = 1;
localparam QSFP2_TEMPERATURE = 'h8a;
localparam QSFP2_TEMPERATURE_SIZE = 2;
localparam QSFP2_VSUPPLY = 'h8c;
localparam QSFP2_VSUPPLY_SIZE = 2;
localparam QSFP2_RXPOWER = 'h8e;
localparam QSFP2_RXPOWER_SIZE = 8;
localparam QSFP2_IDENTIFIER = 'h96;
localparam QSFP2_IDENTIFIER_SIZE = 2;
