module cctrl_marble_top #(
  parameter PILOT_TONE_REFERENCE_DIRECT_OUTPUT_ENABLE = "false"
  ) (
  input              DDR_REF_CLK_P, // 125 MHz
  input              DDR_REF_CLK_N, // 125 MHz (complement)
  //output             VCXO_EN,
  output             PHY_RSTN,

  input  wire        FPGA_TxD,
  output wire        FPGA_RxD,

  input wire         MGT_CLK_1_N, MGT_CLK_1_P,
  input wire         MGT_CLK_2_N, MGT_CLK_2_P,

  input              RGMII_RX_CLK,
  input              RGMII_RX_CTRL,
  input        [3:0] RGMII_RXD,
  output wire        RGMII_TX_CLK,
  output wire        RGMII_TX_CTRL,
  output wire  [3:0] RGMII_TXD,

/*
  Transceiver Assignments (Kintex-7):
  -----------------------------------
    This is copied directly from
      https://controls.als.lbl.gov/alscg/beampositionmonitor/BPM_CC/Documents/HardwareNotes.html

    RX N/P  TX N/P  Tile  MGT           Fiber Pair  QSFP (BMB7) QSFP (Marble)  Desc.
    --------------------------------------------------------------------------------
    C3/C4   B1/B2   X0Y6  MGT2 Bank 116 1:12        1-0         1-1             EVR
    B5/B6   A3/A4   X0Y7  MGT3 Bank 116 2:11        1-1         1-3             BPM CCW
    E3/E4   D1/D2   X0Y5  MGT1 Bank 116 3:10        1-2         1-0             BPM CW
    G3/G4   F1/F2   X0Y4  MGT0 Bank 116 4:9         1-3         1-2             (Unused)
    L3/L4   K1/K2   X0Y2  MGT2 Bank 115 1:12        2-0         2-1             Cell CCW
    J3/J4   H1/H2   X0Y3  MGT3 Bank 115 2:11        2-1         2-3             Cell CW
    N3/N4   M1/M2   X0Y1  MGT1 Bank 115 3:10        2-2         2-0             FOFB power supply chain head (Tx)
    R3/R4   P1/P2   X0Y0  MGT0 Bank 115 4:9         2-3         2-2             FOFB power supply chain tail (Rx)
*/

  input  wire  [2:0] QSFP1_RX_N, QSFP1_RX_P, // [0]->EVR;     [1]->BPM_CCW_GT_RX_rxn; [2]->BPM_CW_GT_RX_rxn
  output wire  [2:1] QSFP1_TX_N, QSFP1_TX_P, // [0]->Unused;  [1]->BPM_CCW; [2]->BPM_CW
  input  wire  [3:0] QSFP2_RX_N, QSFP2_RX_P, // [0]->CELL_CCW_GT_RX_rxn; [1]->CELL_CW_GT_RX_rxn; [2]->fofb(psTx); [3]->fofb(psRx)
  output wire  [3:0] QSFP2_TX_N, QSFP2_TX_P, // [0]->CELL_CCW_GT_TX_txn; [1]->CELL_CW_GT_TX_txn; [2]->fofb(psTx); [3]->fofb(psRx)

  inout TWI_SDA,
  inout TWI_SCL,
  inout TWI_SW_RST,
  // Pinout to match PmodUSBUART (strangely, not Pmod UART standard)
  input PMOD1_0,  // SCRAP ~CTS from USB-UART ~RTS (Unused)
  output PMOD1_1, // SCRAP TxD to USB-UART RxD
  input PMOD1_2,  // SCRAP RxD from USB-UART TxD
  output PMOD1_3, // SCRAP ~RTS to USB-UART ~CTS (Unused)

  output PMOD2_0,
  output PMOD2_1,
  output PMOD2_2,
  output PMOD2_3,
  output PMOD2_4,
  output PMOD2_5,
  output PMOD2_6,
  output PMOD2_7,

  output wire        MARBLE_LD16,
  output wire        MARBLE_LD17
);

wire gtReset = 1'b0;
wire INTLK_RELAY_NO = 1'b0;
wire INTLK_RELAY_CTL;
wire INTLK_RESET_BUTTON_N = 1'b0;

wire FP_LED0_RED, FP_LED0_GRN;  // TODO - Will these exist on marble port?
wire FP_LED1_RED, FP_LED1_GRN;  // TODO - Will these exist on marble port?
wire FP_LED2_RED, FP_LED2_GRN;  // TODO - Will these exist on marble port?
assign PHY_RSTN = 1'b1; // Release the ethernet PHY from reset


//////////////////////////////////////////////////////////////////////////////
// Static outputs

//////////////////////////////////////////////////////////////////////////////
// The clock domains
// Net names starting with 'evr' are in the event receiver clock domain.
// Net names starting with 'aurora' are in the Aurora user clock domain.

wire evrClk;    // Recovered Rx clock from EVR MGT block
wire auroraUserClk; // Generated by Aurora block in 'system' BD

parameter SYSCLK_RATE   = 100_000_000;
parameter FREQ_CLKIN_HZ = 125_000_000;
wire clkIn125;  // Input clock (125 MHz) from U20
wire sysClk;    // 100 MHz sysclk
wire clk200;    // 200 MHz clock
wire ethernetRxClk, ethernetTxClk;
wire ethRefClk125, ethRefClk125Buff;
wire badgerRefClk125, badgerRefClk125d90; // 125 MHz ethernet clock (and 90-deg shifted copy)
wire sysReset_n;

/*
 * 600MHz <= F_VCO <= 1200 MHz
 * F_VCO  = F_CLKIN * CLKFBOUT_MULT_F/DIVCLK_DIVIDE
 * F_OUTx = F_VCO/CLKOUTx_DIVIDE
 *
 * Cell-controller bmb7 port wants 3 output frequencies:
 *   50 MHz, 100 MHz, 200 MHz
 * Ethernet RGMII wants 125 MHz
 * Input is 125MHz
 *
 * Least Common Multiple (LCM) = 1000 MHz
 * F_CLKIN = 125MHz
 *  F_VCO = LCM = 1000 MHz
 *  CLKFBOUT_MULT_F = 8
 *
 * CLKOUT0 = 125 MHz 0deg     => badgerRefClk125
 *  CLKOUT0_DIVIDE = 8
 * CLKOUT1 = 125 MHz 90deg    => badgerRefClk125d90
 *  CLKOUT1_DIVIDE = 8
 * CLKOUT2 = 200 MHz 0deg     => clk200
 *  CLKOUT2_DIVIDE = 5
 * CLKOUT3 = 100 MHz 0deg     => sysClk
 *  CLKOUT3_DIVIDE = 10
 * CLKOUT4 =  50 MHz 0deg     => clk50
 *  CLKOUT4_DIVIDE = 20
 */

IBUFGDS ibufgds_i (
  .O  (clkIn125),
  .I  (DDR_REF_CLK_P),
  .IB (DDR_REF_CLK_N)
);

//////////////////////////////////////////////////////////////////////////////
// General-purpose I/O block
`include "gpioIDX.vh"
wire                    [31:0] GPIO_IN[0:GPIO_IDX_COUNT-1];
wire                    [31:0] GPIO_OUT;
wire      [GPIO_IDX_COUNT-1:0] GPIO_STROBES;
wire [(GPIO_IDX_COUNT*32)-1:0] GPIO_IN_FLATTENED;
genvar i;
generate
for (i = 0 ; i < GPIO_IDX_COUNT ; i = i + 1) begin : gpio_flatten
    assign GPIO_IN_FLATTENED[ (i*32)+31 : (i*32)+0 ] = GPIO_IN[i];
end
endgenerate

//////////////////////////////////////////////////////////////////////////////
// Timekeeping
reg [31:0] secondsSinceBoot, microsecondsSinceBoot;
reg [$clog2(SYSCLK_RATE/1000000)-1:0] microsecondsDivider=SYSCLK_RATE/1000000-1;
reg             [$clog2(1000000)-1:0] secondsDivider = 1000000-1;
reg usTick = 0, sTick = 0;
always @(posedge sysClk) begin
    if (microsecondsDivider == 0) begin
        microsecondsDivider <= SYSCLK_RATE/1000000-1;
        usTick <= 1;
    end
    else begin
        microsecondsDivider <= microsecondsDivider - 1;
        usTick <= 0;
    end
    if (usTick) begin
        microsecondsSinceBoot <= microsecondsSinceBoot + 1;
        if (secondsDivider == 0) begin
            secondsDivider <= 1000000-1;
            sTick <= 1;
        end
        else begin
            secondsDivider <= secondsDivider - 1;
        end
    end
    else begin
        sTick <= 0;
    end
    if (sTick) begin
        secondsSinceBoot <= secondsSinceBoot + 1;
    end
end
assign GPIO_IN[GPIO_IDX_SECONDS]      = secondsSinceBoot;
assign GPIO_IN[GPIO_IDX_MICROSECONDS] = microsecondsSinceBoot;

// Get EVR timestamp to system clock domain
wire [63:0] evrTimestamp, sysTimestamp;
forwardData #(.DATA_WIDTH(64))
  forwardData(.inClk(evrClk),
              .inData(evrTimestamp),
              .outClk(sysClk),
              .outData(sysTimestamp));

wire i2c_run_stat;
wire qsfp_led;
wire qsfp_scl_mon;
wire qsfp_sda_mon;
wire busmux_reset;
wire busmux_reset_i;
IOBUF iobuf_sw_rst(.T(~busmux_reset), .I(1'b0), .O(busmux_reset_i), .IO(TWI_SW_RST));

reg qsfp_freeze=1'b0;
`ifdef QSFP_DEBUG_BUS
//////////////////////////////////////////////////////////////////////////////
// SCRAP Debug Memory Interface

// Bypass hardware flow control
assign PMOD1_3 = 1'b0; // SCRAP ~RTS to USB-UART ~CTS

localparam F_BAUD = 115200;
localparam SCRAP_ADDRESS_WIDTH = 16;
localparam SCRAP_DATA_WIDTH = 8;
wire ext_uart_txd_out;
wire ext_uart_rxd_in = PMOD1_2;
assign PMOD1_1 = ext_uart_txd_out;
wire [SCRAP_ADDRESS_WIDTH-1:0] scrap_addr;
wire [SCRAP_DATA_WIDTH-1:0] scrap_rdata;
wire [SCRAP_DATA_WIDTH-1:0] scrap_wdata;
wire scrap_we;
wire scrap_bus_claim;
wire scrap_bus_claimed = scrap_bus_claim; // SCRAP dev has priority
scrap_dev #(
  .F_CLK_IN(SYSCLK_RATE),
  .F_BAUD(F_BAUD),
  .ADDRESS_WIDTH(SCRAP_ADDRESS_WIDTH),
  .DATA_WIDTH(SCRAP_DATA_WIDTH),
  .LATCH_CYCLES(2)
) scrap_dev_inst (
  .clk(sysClk),
  .rst(1'b0),
  // PHY interface
  .uart_rxd(ext_uart_rxd_in),   // input
  .uart_txd(ext_uart_txd_out),  // output
  // Memory interface
  .addr(scrap_addr),    // output [ADDRESS_WIDTH-1:0]
  .rdata(scrap_rdata),  // input [DATA_WIDTH-1:0]
  .wdata(scrap_wdata),  // output [DATA_WIDTH-1:0]
  .we(scrap_we),
  .op(),
  // Shared bus
  .bus_claim(scrap_bus_claim),  // output
  .bus_claimed(scrap_bus_claimed),  // input
  // Status
  .error_count()
);

wire [7:0] qsfp_lb_dout;
reg qsfp_run_cmd;
reg [7:0] scrap_rdata_hi;
initial begin
  qsfp_run_cmd = 1'b1;
  qsfp_freeze = 1'b0;
  scrap_rdata_hi = 0;
end
// Memory map
wire qsfp_we = scrap_addr[12] ? 1'b0 : scrap_we;
assign scrap_rdata = scrap_addr[12] ? scrap_rdata_hi : qsfp_lb_dout;

always @(posedge sysClk) begin
  if (scrap_we) begin
    case (scrap_addr)
      'h1000 : {qsfp_freeze, qsfp_run_cmd} <= scrap_wdata[1:0];
    endcase
  end
  case (scrap_addr)
    'h1000 : scrap_rdata_hi <= {5'h0, busmux_reset_i, qsfp_buffer_freeze, i2c_run_stat};
    default: scrap_rdata_hi <= 8'h00;
  endcase
end

assign PMOD2_0 = qsfp_run_cmd;
assign PMOD2_1 = i2c_run_stat;
assign PMOD2_2 = scrap_we;
assign PMOD2_3 = qsfp_led;
assign PMOD2_4 = qsfp_scl_mon;
assign PMOD2_5 = qsfp_sda_mon;
assign PMOD2_6 = i2c_updated;
assign PMOD2_7 = 1'b0;
`else
assign PMOD2_0 = 1'b0;
assign PMOD2_1 = 1'b0;
assign PMOD2_2 = 1'b0;
assign PMOD2_3 = 1'b0;
assign PMOD2_4 = 1'b0;
assign PMOD2_5 = 1'b0;
assign PMOD2_6 = 1'b0;
assign PMOD2_7 = 1'b0;
`endif

//////////////////////////////////////////////////////////////////////////////
// QSFP monitoring
parameter QSFP_COUNT = 2;
reg [$clog2(QSFP_COUNT)+7:0] qsfpReadAddress;
reg i2c_buffer_freeze;
initial begin
  qsfpReadAddress = 0;
  i2c_buffer_freeze = 1'b0;
end
wire [7:0] qsfpReadData;
wire i2c_updated;
assign GPIO_IN[GPIO_IDX_QSFP_IIC] = {{22{1'b0}}, i2c_updated, i2c_run_stat, qsfpReadData};
always @(posedge sysClk) begin
    if (GPIO_STROBES[GPIO_IDX_QSFP_IIC]) begin
        qsfpReadAddress <= GPIO_OUT[$clog2(QSFP_COUNT)+7:0];
        i2c_buffer_freeze <= GPIO_OUT[16];
    end
end

wire qsfp_buffer_freeze = qsfp_freeze | i2c_buffer_freeze;
qsfpMarble #(
  .QSFP_COUNT(QSFP_COUNT),
  .CLOCK_RATE(SYSCLK_RATE),
  .BIT_RATE(100000)
  ) qsfpMarble_i (
  .clk(sysClk), // input
  .readAddress(qsfpReadAddress), // input [$clog2(QSFP_COUNT)+7:0]
  .readData(qsfpReadData), // output [7:0]
  .freeze(qsfp_buffer_freeze), // input
  .run_stat(i2c_run_stat), // output
  .updated(i2c_updated), // output
  .SCL(TWI_SCL), // inout
  .SDA(TWI_SDA), // inout
  .scl_mon(qsfp_scl_mon),
  .sda_mon(qsfp_sda_mon),
`ifdef QSFP_DEBUG_BUS
  .bus_claim(scrap_bus_claim),
  .lb_addr(scrap_addr[11:0]), // input [11:0]
  .lb_din(scrap_wdata),
  .lb_dout(qsfp_lb_dout),
  .lb_write(qsfp_we),
  .run_cmd(qsfp_run_cmd),
`endif
  .led(qsfp_led),
  .busmux_reset(busmux_reset)
);

/////////////////////////////////////////////////////////////////////////////
// Event receiver
wire [7:0] evrTriggerBus, evrDataBus;
wire evrFAmarker, evrIsSynchronized, evrHeartbeatPresent;
reg sysFAenable = 0, evrFAenable_m, evrFAenable;
evrSync evrSync(.clk(evrClk),
                .triggerIn(evrTriggerBus[0]),
                .FAenable(evrFAenable),
                .FAmarker(evrFAmarker),
                .isSynchronized(evrIsSynchronized),
                .triggered(evrHeartbeatPresent));
assign GPIO_IN[GPIO_IDX_EVENT_STATUS] = { 29'b0,
                                          evrRxLocked,
                                          evrIsSynchronized,
                                          evrHeartbeatPresent };
always @(posedge evrClk) begin
    evrFAenable_m <= sysFAenable;
    evrFAenable   <= evrFAenable_m;
end
reg auroraFAmarker_m, auroraFAmarker, auroraFAmarker_d, auroraFAstrobe;
always @(posedge auroraUserClk) begin
    auroraFAmarker_m <= evrFAmarker;
    auroraFAmarker   <= auroraFAmarker_m;
    auroraFAmarker_d <= auroraFAmarker;
    auroraFAstrobe <= (auroraFAmarker && !auroraFAmarker_d);
end
reg sysFAmarker_m, sysFAmarker, sysFAmarker_d, sysFAstrobe;
always @(posedge sysClk) begin
    sysFAmarker_m <= evrFAmarker;
    sysFAmarker   <= sysFAmarker_m;
    sysFAmarker_d <= sysFAmarker;
    sysFAstrobe <= (sysFAmarker && !sysFAmarker_d);
end

//////////////////////////////////////////////////////////////////////////////
// BPM and cell readout
wire pll_not_locked_out, gt0_qplllock_out, gt0_qpllrefclklost_out, gtxResetOut;
reg sysGTXreset = 1, sysAuroraReset = 1, auroraReset_m = 1, auroraReset = 1;
always @(posedge sysClk) begin
    if (GPIO_STROBES[GPIO_IDX_AURORA_CSR]) begin
        sysGTXreset    <= GPIO_OUT[0];
        sysAuroraReset <= GPIO_OUT[1];
        sysFAenable    <= GPIO_OUT[2];
    end
end
always @(posedge auroraUserClk) begin
    auroraReset_m <= sysAuroraReset;
    auroraReset   <= auroraReset_m;
end
assign GPIO_IN[GPIO_IDX_AURORA_CSR] = { 8'b0,
     CELL_CW_AuroraCoreStatus_hard_err, CELL_CCW_AuroraCoreStatus_hard_err,
     BPM_CW_AuroraCoreStatus_hard_err, BPM_CCW_AuroraCoreStatus_hard_err,
     CELL_CW_AuroraCoreStatus_soft_err, CELL_CCW_AuroraCoreStatus_soft_err,
     BPM_CW_AuroraCoreStatus_soft_err, BPM_CCW_AuroraCoreStatus_soft_err,
     CELL_CW_AuroraCoreStatus_channel_up, CELL_CCW_AuroraCoreStatus_channel_up,
     BPM_CW_AuroraCoreStatus_channel_up, BPM_CCW_AuroraCoreStatus_channel_up,
     pll_not_locked_out, gt0_qplllock_out, gt0_qpllrefclklost_out, gtxResetOut,
     5'b0, sysFAenable, sysAuroraReset, sysGTXreset };

/////////////////////////////////////////////////////////////////////////////
// Event receiver GTX
localparam EVR_DEBUG = "false";
wire        evr_mgt_drp_den, evr_mgt_drp_drdy, evr_mgt_drp_dwe;
wire [15:0] evr_mgt_drp_di, evr_mgt_drp_do;
wire  [8:0] evr_mgt_drp_daddr;
(* mark_debug=EVR_DEBUG *) wire  [1:0] evr_mgt_chariscomma, evr_mgt_charisk;
(* mark_debug=EVR_DEBUG *) wire  [1:0] evr_notintable;
(* mark_debug=EVR_DEBUG *) wire [15:0] evr_mgt_par_data;
(* mark_debug=EVR_DEBUG *) wire        evr_mgt_reset_done;

evr_mgt_top #(.COMMA_IS_LSB_FORCE(1)) evr_mgt_top_i (
         .reset(gtReset),
         .ref_clk(ethRefClk125),  // Comes from bank 115
         .drp_clk(sysClk),
         .drp_den(evr_mgt_drp_den),
         .drp_dwe(evr_mgt_drp_dwe),
         .drp_daddr(evr_mgt_drp_daddr),
         .drp_di(evr_mgt_drp_di),
         .drp_drdy(evr_mgt_drp_drdy),
         .drp_do(evr_mgt_drp_do),
         .rx_in_n(QSFP1_RX_N[0]), // Bank 116!
         .rx_in_p(QSFP1_RX_P[0]), // Bank 116!
         .rec_clk_out(evrClk),
         .rx_par_data_out(evr_mgt_par_data),
         .chariscomma(evr_mgt_chariscomma),
         .notintable(evr_notintable),
         .charisk(evr_mgt_charisk),
         .reset_done(evr_mgt_reset_done));

// Announce that receiver clock is locked only when all
// characters have been valid 8b/10b codes for a while.
(* mark_debug = EVR_DEBUG *) reg       evrRxLocked = 0;
                             reg [3:0] evrGoodCount = 0;
always @(posedge evrClk) begin
    if (|evr_notintable) begin
        evrRxLocked <= 0;
        evrGoodCount <= 0;
    end
    else if (evrGoodCount == 15) begin
        evrRxLocked <= 1;
    end
    else begin
        evrGoodCount <= evrGoodCount + 1;
    end
end

//////////////////////////////////////////////////////////////////////////////
// Event stream logger
evrLogger #(.ADDR_WIDTH(8))
  evrLogger (
    .sysClk(sysClk),
    .sysCsrStrobe(GPIO_STROBES[GPIO_IDX_EVENT_LOG_CSR]),
    .sysGpioOut(GPIO_OUT),
    .sysCsr(GPIO_IN[GPIO_IDX_EVENT_LOG_CSR]),
    .sysDataTicks(GPIO_IN[GPIO_IDX_EVENT_LOG_TICKS]),
    .evrClk(evrClk),
    .evrTVALID(!evr_mgt_charisk[0]),
    .evrTDATA(evr_mgt_par_data[7:0]));

//////////////////////////////////////////////////////////////////////////////
// Aurora streams

// BPM CCW link
wire        BPM_CCW_AXI_STREAM_RX_tlast, BPM_CCW_AXI_STREAM_RX_tvalid;
wire [31:0] BPM_CCW_AXI_STREAM_RX_tdata;
wire        BPM_CCW_AuroraCoreStatus_channel_up;
wire        BPM_CCW_AuroraCoreStatus_crc_pass_fail;
wire        BPM_CCW_AuroraCoreStatus_crc_valid;
wire        BPM_CCW_AuroraCoreStatus_frame_err;
wire        BPM_CCW_AuroraCoreStatus_hard_err;
wire        BPM_CCW_AuroraCoreStatus_lane_up;
wire        BPM_CCW_AuroraCoreStatus_rx_resetdone_out;
wire        BPM_CCW_AuroraCoreStatus_soft_err;
wire        BPM_CCW_AuroraCoreStatus_tx_lock;
wire        BPM_CCW_AuroraCoreStatus_tx_resetdone_out;

// BPM CW link
wire        BPM_CW_AXI_STREAM_RX_tlast, BPM_CW_AXI_STREAM_RX_tvalid;
wire [31:0] BPM_CW_AXI_STREAM_RX_tdata;
wire        BPM_CW_AuroraCoreStatus_channel_up;
wire        BPM_CW_AuroraCoreStatus_crc_pass_fail;
wire        BPM_CW_AuroraCoreStatus_crc_valid;
wire        BPM_CW_AuroraCoreStatus_frame_err;
wire        BPM_CW_AuroraCoreStatus_hard_err;
wire        BPM_CW_AuroraCoreStatus_lane_up;
wire        BPM_CW_AuroraCoreStatus_rx_resetdone_out;
wire        BPM_CW_AuroraCoreStatus_soft_err;
wire        BPM_CW_AuroraCoreStatus_tx_lock;
wire        BPM_CW_AuroraCoreStatus_tx_resetdone_out;

// Cell CCW link
localparam CELL_AXI_DEBUG = "false";
(* mark_debug = CELL_AXI_DEBUG *) wire        CELL_CCW_AXI_STREAM_TX_tvalid;
(* mark_debug = CELL_AXI_DEBUG *) wire        CELL_CCW_AXI_STREAM_TX_tready;
(* mark_debug = CELL_AXI_DEBUG *) wire        CELL_CCW_AXI_STREAM_TX_tlast;
(* mark_debug = CELL_AXI_DEBUG *) wire [31:0] CELL_CCW_AXI_STREAM_TX_tdata;
(* mark_debug = CELL_AXI_DEBUG *) wire        CELL_CCW_AXI_STREAM_RX_tvalid;
(* mark_debug = CELL_AXI_DEBUG *) wire        CELL_CCW_AXI_STREAM_RX_tlast;
(* mark_debug = CELL_AXI_DEBUG *) wire [31:0] CELL_CCW_AXI_STREAM_RX_tdata;
wire        CELL_CCW_AuroraCoreStatus_channel_up;
wire        CELL_CCW_AuroraCoreStatus_crc_pass_fail;
wire        CELL_CCW_AuroraCoreStatus_crc_valid;
wire        CELL_CCW_AuroraCoreStatus_frame_err;
wire        CELL_CCW_AuroraCoreStatus_hard_err;
wire        CELL_CCW_AuroraCoreStatus_lane_up;
wire        CELL_CCW_AuroraCoreStatus_rx_resetdone_out;
wire        CELL_CCW_AuroraCoreStatus_soft_err;
wire        CELL_CCW_AuroraCoreStatus_tx_lock;
wire        CELL_CCW_AuroraCoreStatus_tx_resetdone_out;

// Cell CW link
(* mark_debug = CELL_AXI_DEBUG *) wire        CELL_CW_AXI_STREAM_TX_tvalid;
(* mark_debug = CELL_AXI_DEBUG *) wire        CELL_CW_AXI_STREAM_TX_tready;
(* mark_debug = CELL_AXI_DEBUG *) wire        CELL_CW_AXI_STREAM_TX_tlast;
(* mark_debug = CELL_AXI_DEBUG *) wire [31:0] CELL_CW_AXI_STREAM_TX_tdata;
(* mark_debug = CELL_AXI_DEBUG *) wire        CELL_CW_AXI_STREAM_RX_tvalid;
(* mark_debug = CELL_AXI_DEBUG *) wire        CELL_CW_AXI_STREAM_RX_tlast;
(* mark_debug = CELL_AXI_DEBUG *) wire [31:0] CELL_CW_AXI_STREAM_RX_tdata;
wire        CELL_CW_AuroraCoreStatus_channel_up;
wire        CELL_CW_AuroraCoreStatus_crc_pass_fail;
wire        CELL_CW_AuroraCoreStatus_crc_valid;
wire        CELL_CW_AuroraCoreStatus_frame_err;
wire        CELL_CW_AuroraCoreStatus_hard_err;
wire        CELL_CW_AuroraCoreStatus_lane_up;
wire        CELL_CW_AuroraCoreStatus_rx_resetdone_out;
wire        CELL_CW_AuroraCoreStatus_soft_err;
wire        CELL_CW_AuroraCoreStatus_tx_lock;
wire        CELL_CW_AuroraCoreStatus_tx_resetdone_out;

//////////////////////////////////////////////////////////////////////////////
// Read and coalesce data from BPM links
wire [31:0] localBPMs_tdata;
wire        localBPMs_tvalid, localBPMs_tlast;
wire  [1:0] bpmCCWstatusCode,    bpmCWstatusCode;
wire        bpmCCWstatusStrobe,  bpmCWstatusStrobe;
wire  [2:0] sysCellStatusCode;
wire        sysCellStatusStrobe;

wire [111:0] localBPMvalues;      // Aurora user clock domain
wire         localBPMvaluesVALID; // Aurora user clock domain

wire [31:0] BRAM_BPM_SETPOINTS_WDATA;
wire [15:0] BRAM_BPM_SETPOINTS_ADDR;
wire        BRAM_BPM_SETPOINTS_WENABLE;
wire [31:0] BRAM_BPM_SETPOINTS_RDATA;

reg localFOFBcontrol = 0;
wire fofbEnabled;
always @(posedge sysClk) begin
    if (GPIO_STROBES[GPIO_IDX_FOFB_CSR]) localFOFBcontrol <= GPIO_OUT[0];
end
assign GPIO_IN[GPIO_IDX_FOFB_CSR] = {{29{1'b0}},
                               fofbEnabled, 1'b0, localFOFBcontrol};

readBPMlinks #(.faStrobeDebug("false"),
               .bpmSetpointDebug("false"),
               .ccwInDebug("false"),
               .cwInDebug("false"),
               .mergedDebug("false"),
               .outDebug("false"),
               .stateDebug("false"))
  readBPMlinks (
         .sysClk(sysClk),
         .sysCsrStrobe(GPIO_STROBES[GPIO_IDX_BPMLINKS_CSR]),
         .GPIO_OUT(GPIO_OUT),
         .sysCsr(GPIO_IN[GPIO_IDX_BPMLINKS_CSR]),
         .sysAdditionalStatus(GPIO_IN[GPIO_IDX_BPMLINKS_EXTRA_STATUS]),
         .sysRxBitmap(GPIO_IN[GPIO_IDX_BPM_RX_BITMAP]),
         .sysLocalFOFBenabled(localFOFBcontrol),
         .sysSetpointWriteData(BRAM_BPM_SETPOINTS_WDATA),
         .sysSetpointAddress(BRAM_BPM_SETPOINTS_ADDR),
         .sysSetpointWriteEnable(BRAM_BPM_SETPOINTS_WENABLE),
         .sysSetpointReadData(BRAM_BPM_SETPOINTS_RDATA),
         .auroraUserClk(auroraUserClk),
         .auroraFAstrobe(auroraFAstrobe),
         .BPM_CCW_AXI_STREAM_RX_tdata(BPM_CCW_AXI_STREAM_RX_tdata),
         .BPM_CCW_AXI_STREAM_RX_tvalid(BPM_CCW_AXI_STREAM_RX_tvalid),
         .BPM_CCW_AXI_STREAM_RX_tlast(BPM_CCW_AXI_STREAM_RX_tlast),
         .BPM_CCW_AXI_STREAM_RX_CRC_pass(BPM_CCW_AuroraCoreStatus_crc_pass_fail),
         .BPM_CCW_AXI_STREAM_RX_CRC_valid(BPM_CCW_AuroraCoreStatus_crc_valid),
         .CCWstatusStrobe(bpmCCWstatusStrobe),
         .CCWstatusCode(bpmCCWstatusCode),
         .BPM_CW_AXI_STREAM_RX_tdata(BPM_CW_AXI_STREAM_RX_tdata),
         .BPM_CW_AXI_STREAM_RX_tvalid(BPM_CW_AXI_STREAM_RX_tvalid),
         .BPM_CW_AXI_STREAM_RX_tlast(BPM_CW_AXI_STREAM_RX_tlast),
         .BPM_CW_AXI_STREAM_RX_CRC_pass(BPM_CW_AuroraCoreStatus_crc_pass_fail),
         .BPM_CW_AXI_STREAM_RX_CRC_valid(BPM_CW_AuroraCoreStatus_crc_valid),
         .CWstatusStrobe(bpmCWstatusStrobe),
         .CWstatusCode(bpmCWstatusCode),
         .mergedLinkTDATA(localBPMvalues),
         .mergedLinkTVALID(localBPMvaluesVALID),
         .localBPMs_tdata(localBPMs_tdata),
         .localBPMs_tvalid(localBPMs_tvalid),
         .localBPMs_tlast(localBPMs_tlast));

//////////////////////////////////////////////////////////////////////////////
// Forward incoming and local streams to next cell
// Pick up CSR values from fofbReadLinks since we don't have any CSR
wire auCCWcellInhibit, auCWcellInhibit;
wire auCCWcellStreamValid = CELL_CCW_AXI_STREAM_RX_tvalid && !auCCWcellInhibit;
wire auCWcellStreamValid  = CELL_CW_AXI_STREAM_RX_tvalid  && !auCWcellInhibit;
forwardCellLink #(.dbg("false")) forwardCCWcell (
       .auroraUserClk(auroraUserClk),
       .auroraFAstrobe(auroraFAstrobe),
       .cellLinkRxTVALID(auCCWcellStreamValid),
       .cellLinkRxTLAST(CELL_CCW_AXI_STREAM_RX_tlast),
       .cellLinkRxTDATA(CELL_CCW_AXI_STREAM_RX_tdata),
       .cellLinkRxCRCvalid(CELL_CCW_AuroraCoreStatus_crc_valid),
       .cellLinkRxCRCpass(CELL_CCW_AuroraCoreStatus_crc_pass_fail),
       .localRxTVALID(localBPMs_tvalid),
       .localRxTLAST(localBPMs_tlast),
       .localRxTDATA(localBPMs_tdata),
       .cellLinkTxTVALID(CELL_CW_AXI_STREAM_TX_tvalid),
       .cellLinkTxTLAST(CELL_CW_AXI_STREAM_TX_tlast),
       .cellLinkTxTDATA(CELL_CW_AXI_STREAM_TX_tdata));
forwardCellLink #(.dbg("false")) forwardCWcell (
       .auroraUserClk(auroraUserClk),
       .auroraFAstrobe(auroraFAstrobe),
       .cellLinkRxTVALID(auCWcellStreamValid),
       .cellLinkRxTLAST(CELL_CW_AXI_STREAM_RX_tlast),
       .cellLinkRxTDATA(CELL_CW_AXI_STREAM_RX_tdata),
       .cellLinkRxCRCvalid(CELL_CW_AuroraCoreStatus_crc_valid),
       .cellLinkRxCRCpass(CELL_CW_AuroraCoreStatus_crc_pass_fail),
       .localRxTVALID(localBPMs_tvalid),
       .localRxTLAST(localBPMs_tlast),
       .localRxTDATA(localBPMs_tdata),
       .cellLinkTxTVALID(CELL_CCW_AXI_STREAM_TX_tvalid),
       .cellLinkTxTLAST(CELL_CCW_AXI_STREAM_TX_tlast),
       .cellLinkTxTDATA(CELL_CCW_AXI_STREAM_TX_tdata));

//////////////////////////////////////////////////////////////////////////////
// Gather data from outgoing streams and make available to fast orbit feedback
wire        sysTimeoutStrobe;
wire [31:0] fofbReadoutCSR, fofbDSPreadoutS, fofbDSPreadoutY, fofbDSPreadoutX;
wire [GPIO_FOFB_MATRIX_ADDR_WIDTH-1:0] fofbDSPreadoutAddress;
assign GPIO_IN[GPIO_IDX_CELL_COMM_CSR] = fofbReadoutCSR;
fofbReadLinks #(.SYSCLK_RATE(SYSCLK_RATE),
                .FOFB_INDEX_WIDTH(GPIO_FOFB_MATRIX_ADDR_WIDTH),
                .FAstrobeDebug("false"),
                .statusDebug("false"),
                .rawDataDebug("false"),
                .ccwLinkDebug("false"),
                .cwLinkDebug("false"),
                .cellCountDebug("false"),
                .dspReadoutDebug("false"))
  fofbReadLinks (
       .sysClk(sysClk),
       .csrStrobe(GPIO_STROBES[GPIO_IDX_CELL_COMM_CSR]),
       .GPIO_OUT(GPIO_OUT),
       .csr(fofbReadoutCSR),
       .rxBitmap(GPIO_IN[GPIO_IDX_CELL_RX_BITMAP]),
       .fofbEnableBitmap(GPIO_IN[GPIO_IDX_FOFB_ENABLE_BITMAP]),
       .fofbEnabled(fofbEnabled),

       .FAstrobe(sysFAstrobe),
       .auReset(auroraReset),
       .sysStatusStrobe(sysCellStatusStrobe),
       .sysStatusCode(sysCellStatusCode),
       .sysTimeoutStrobe(sysTimeoutStrobe),

       .fofbDSPreadoutAddress(fofbDSPreadoutAddress),
       .fofbDSPreadoutX(fofbDSPreadoutX),
       .fofbDSPreadoutY(fofbDSPreadoutY),
       .fofbDSPreadoutS(fofbDSPreadoutS),

       .uBreadoutStrobe(GPIO_STROBES[GPIO_IDX_BPM_READOUT_X]),
       .uBreadoutX(GPIO_IN[GPIO_IDX_BPM_READOUT_X]),
       .uBreadoutY(GPIO_IN[GPIO_IDX_BPM_READOUT_Y]),
       .uBreadoutS(GPIO_IN[GPIO_IDX_BPM_READOUT_S]),

       .auClk(auroraUserClk),
       .auFAstrobe(auroraFAstrobe),
       .auCCWcellInhibit(auCCWcellInhibit),
       .auCWcellInhibit(auCWcellInhibit),

       .auCellCCWlinkTVALID(CELL_CCW_AXI_STREAM_TX_tvalid),
       .auCellCCWlinkTLAST(CELL_CCW_AXI_STREAM_TX_tlast),
       .auCellCCWlinkTDATA(CELL_CCW_AXI_STREAM_TX_tdata),

       .auCellCWlinkTVALID(CELL_CW_AXI_STREAM_TX_tvalid),
       .auCellCWlinkTLAST(CELL_CW_AXI_STREAM_TX_tlast),
       .auCellCWlinkTDATA(CELL_CW_AXI_STREAM_TX_tdata));

//////////////////////////////////////////////////////////////////////////////
// Keep link reception statistics
linkStatistics #(.dbg("false")) linkStatistics (
         .auroraUserClk(auroraUserClk),
         .bpmCCWstatusStrobe(bpmCCWstatusStrobe),
         .bpmCCWstatusCode  (bpmCCWstatusCode),
         .bpmCWstatusStrobe (bpmCWstatusStrobe),
         .bpmCWstatusCode   (bpmCWstatusCode),
         .sysClk(sysClk),
         .sysStatusStrobe (sysCellStatusStrobe),
         .sysStatusCode   (sysCellStatusCode),
         .sysTimeoutStrobe(sysTimeoutStrobe),
         .sysCsrStrobe(GPIO_STROBES[GPIO_IDX_LINK_STATISTICS_CSR]),
         .GPIO_OUT(GPIO_OUT),
         .sysValue(GPIO_IN[GPIO_IDX_LINK_STATISTICS_CSR]));

//////////////////////////////////////////////////////////////////////////////
// Compute power supply settings
wire        FOFB_SETPOINT_AXIS_TVALID;
wire        FOFB_SETPOINT_AXIS_TLAST;
wire [31:0] FOFB_SETPOINT_AXIS_TDATA;
fofbDSP #(.RESULT_COUNT(GPIO_CHANNEL_COUNT),
          .FOFB_MATRIX_ADDR_WIDTH(GPIO_FOFB_MATRIX_ADDR_WIDTH),
          .MATMUL_DEBUG("false"),
          .FIR_DEBUG("false"),
          .TX_AXIS_DEBUG("false"))
  fofbDSP (
    .clk(sysClk),
    .csrStrobe(GPIO_STROBES[GPIO_IDX_DSP_CSR]),
    .GPIO_OUT(GPIO_OUT),
    .firStatus(GPIO_IN[GPIO_IDX_DSP_CSR]),
    .fofbReadoutCSR(fofbReadoutCSR),
    .fofbEnabled(fofbEnabled),
    .fofbDSPreadoutAddress(fofbDSPreadoutAddress),
    .fofbDSPreadoutX(fofbDSPreadoutX),
    .fofbDSPreadoutY(fofbDSPreadoutY),
    .fofbDSPreadoutS(fofbDSPreadoutS),
    .SETPOINT_TVALID(FOFB_SETPOINT_AXIS_TVALID),
    .SETPOINT_TLAST(FOFB_SETPOINT_AXIS_TLAST),
    .SETPOINT_TDATA(FOFB_SETPOINT_AXIS_TDATA));

//////////////////////////////////////////////////////////////////////////////
// Provide CPU read access to power supply setpoints
psSetpointMonitor #(.SETPOINT_COUNT(GPIO_CHANNEL_COUNT),
                    .DEBUG("false"))
  psSetpointMonitor (
    .clk(sysClk),
    .FOFB_SETPOINT_AXIS_TVALID(FOFB_SETPOINT_AXIS_TVALID),
    .FOFB_SETPOINT_AXIS_TLAST(FOFB_SETPOINT_AXIS_TLAST),
    .FOFB_SETPOINT_AXIS_TDATA(FOFB_SETPOINT_AXIS_TDATA),
    .addressStrobe(GPIO_STROBES[GPIO_IDX_FOFB_PS_SETPOINT]),
    .GPIO_OUT(GPIO_OUT),
    .psSetpoint(GPIO_IN[GPIO_IDX_FOFB_PS_SETPOINT]),
    .status(GPIO_IN[GPIO_IDX_FOFB_PS_SETPOINT_STATUS]));

//////////////////////////////////////////////////////////////////////////////
// Arbitrary Waveform Generator
wire [31:0] AWG_AXIS_TDATA;
wire        AWG_AXIS_TVALID, AWG_AXIS_TLAST;
wire        AWGrequest, AWGenabled;

psAWG #(.SETPOINT_COUNT(GPIO_CHANNEL_COUNT),
        .DATA_WIDTH(32),
        .ADDR_WIDTH($clog2(GPIO_AWG_CAPACITY)),
        .SYSCLK_RATE(SYSCLK_RATE),
        .DEBUG("false"))
  psAWG (.sysClk(sysClk),
         .csrStrobe(GPIO_STROBES[GPIO_IDX_AWG_CSR]),
         .addrStrobe(GPIO_STROBES[GPIO_IDX_AWG_ADDRESS]),
         .dataStrobe(GPIO_STROBES[GPIO_IDX_AWG_DATA]),
         .GPIO_OUT(GPIO_OUT),
         .status(GPIO_IN[GPIO_IDX_AWG_CSR]),
         .evrTrigger(evrTriggerBus[2]),
         .sysFAstrobe(sysFAstrobe),
         .AWGrequest(AWGrequest),
         .AWGenabled(AWGenabled),
         .awgTDATA(AWG_AXIS_TDATA),
         .awgTVALID(AWG_AXIS_TVALID),
         .awgTLAST(AWG_AXIS_TLAST));

//////////////////////////////////////////////////////////////////////////////
// Multiplex fast feedback and arbitrary waveform streams
wire [31:0] PS_SETPOINT_AXIS_TDATA;
wire        PS_SETPOINT_AXIS_TVALID, PS_SETPOINT_AXIS_TLAST;
wire [31:0] PS_READBACK_AXIS_TDATA;
wire  [7:0] PS_READBACK_AXIS_TUSER;
wire        PS_READBACK_AXIS_TVALID;

psMUX #(.DEBUG("false"),
        .AXI_WIDTH(32))
  psMUX (.clk(sysClk),
         .AWGrequest(AWGrequest),
         .AWGenabled(AWGenabled),
         .fofbTDATA(FOFB_SETPOINT_AXIS_TDATA),
         .fofbTVALID(FOFB_SETPOINT_AXIS_TVALID),
         .fofbTLAST(FOFB_SETPOINT_AXIS_TLAST),
         .awgTDATA(AWG_AXIS_TDATA),
         .awgTVALID(AWG_AXIS_TVALID),
         .awgTLAST(AWG_AXIS_TLAST),
         .psTDATA(PS_SETPOINT_AXIS_TDATA),
         .psTVALID(PS_SETPOINT_AXIS_TVALID),
         .psTLAST(PS_SETPOINT_AXIS_TLAST));

//////////////////////////////////////////////////////////////////////////////
// Ethernet in fabric connection to fast orbit feedback power supplies
// Destination MAC address is as specified in RFC 1112 and RFC 7042:
//               01:00:5E followed by low 23 bits of IPv4 multicast address.
//               IPv4 multicast address is that of the current FastPS firmware:
//                                                                   224.0.2.22.
wire [9:0] pcs_pma_shared;
wire [63:0] ethNonce;
assign  ethRefClk125 = pcs_pma_shared[9];
assign  ethRefClk125Buff = pcs_pma_shared[8];
fofbEthernet #(
    .MAX_CORRECTOR_COUNT(GPIO_CHANNEL_COUNT),
    .PCS_PMA_SHARED_LOGIC_IN_CORE("true"),
    .SRC_IP_ADDRESS({8'd192, 8'd168, 8'd30, 8'd251}),
    .SRC_MAC_ADDRESS({8'h2A,8'h4C,8'h42,8'h4E,8'h4C,8'h32}),
    .DST_MAC_ADDRESS({8'h01, 8'h00, 8'h5E, 8'd0, 8'd2, 8'd22}),
    .DST_IP_ADDRESS(              {8'd224, 8'd0, 8'd2, 8'd22}),
    .TX_DEBUG("false"),
    .RX_DEBUG("false"))
  psTx (
    .sysClk(sysClk),
    .sysGpioOut(GPIO_OUT),
    .sysCsrStrobe(GPIO_STROBES[GPIO_IDX_ETHERNET0_CSR]),
    .sysCsr(GPIO_IN[GPIO_IDX_ETHERNET0_CSR]),
    .sysTx_S_AXIS_TDATA(PS_SETPOINT_AXIS_TDATA),
    .sysTx_S_AXIS_TVALID(PS_SETPOINT_AXIS_TVALID),
    .sysTx_S_AXIS_TLAST(PS_SETPOINT_AXIS_TLAST),
    .pcs_pma_shared(pcs_pma_shared),
    .ethNonce(ethNonce),
    .clk200(clk200),
    .ETH_REF_N(MGT_CLK_2_N),
    .ETH_REF_P(MGT_CLK_2_P),
    .ETH_RX_N(QSFP2_RX_N[2]), // R3  MGT_RX_4_N  MGT_RX_4_QSFP_N   QSFP2_RX_3_N Bank 115
    .ETH_RX_P(QSFP2_RX_P[2]), // R4  MGT_RX_4_P  MGT_RX_4_QSFP_P   QSFP2_RX_3_P Bank 115
    .ETH_TX_N(QSFP2_TX_N[2]), // P1  MGT_TX_4_N  MGT_TX_4_QSFP_N   QSFP2_TX_3_N Bank 115
    .ETH_TX_P(QSFP2_TX_P[2]));// P2  MGT_TX_4_P  MGT_TX_4_QSFP_P   QSFP2_TX_3_P Bank 115

fofbEthernet #(
    .MAX_CORRECTOR_COUNT(GPIO_CHANNEL_COUNT),
    .PCS_PMA_SHARED_LOGIC_IN_CORE("false"),
    .SRC_IP_ADDRESS({8'd192, 8'd168, 8'd30, 8'd250}),
    .SRC_MAC_ADDRESS({8'h2A,8'h4C,8'h42,8'h4E,8'h4C,8'h33}),
    .DST_IP_ADDRESS({8'd255, 8'd255, 8'd255, 8'd255}),
    .DST_MAC_ADDRESS({8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF}),
    .TX_DEBUG("false"),
    .RX_DEBUG("false"))
  psRx (
    .sysClk(sysClk),
    .sysGpioOut(GPIO_OUT),
    .sysCsrStrobe(GPIO_STROBES[GPIO_IDX_ETHERNET1_CSR]),
    .sysCsr(GPIO_IN[GPIO_IDX_ETHERNET1_CSR]),
    .sysTx_S_AXIS_TDATA(32'h0),
    .sysTx_S_AXIS_TVALID(1'b0),
    .sysTx_S_AXIS_TLAST(1'b0),
    .sysRx_M_AXIS_TDATA(PS_READBACK_AXIS_TDATA),
    .sysRx_M_AXIS_TUSER(PS_READBACK_AXIS_TUSER),
    .sysRx_M_AXIS_TVALID(PS_READBACK_AXIS_TVALID),
    .pcs_pma_shared(pcs_pma_shared),
    .ethNonce(ethNonce),
    .clk200(clk200),
    .ETH_REF_N(1'b0),  // NOTE! UNUSED when PCS_PMA_SHARED_LOGIC_IN_CORE == "false"
    .ETH_REF_P(1'b0),  // NOTE! UNUSED when PCS_PMA_SHARED_LOGIC_IN_CORE == "false"
    .ETH_RX_N(QSFP2_RX_N[3]), // J3  MGT_RX_7_N  MGT_RX_7_QSFP_N   QSFP2_RX_4_N Bank 115
    .ETH_RX_P(QSFP2_RX_P[3]), // J4  MGT_RX_7_P  MGT_RX_7_QSFP_P   QSFP2_RX_4_P Bank 115
    .ETH_TX_N(QSFP2_TX_N[3]), // H1  MGT_TX_7_N  MGT_TX_7_QSFP_N   QSFP2_TX_4_N Bank 115
    .ETH_TX_P(QSFP2_TX_P[3]));// H2  MGT_TX_7_P  MGT_TX_7_QSFP_P   QSFP2_TX_4_P Bank 115

//////////////////////////////////////////////////////////////////////////////
// Fast orbit feedback waveform recorder
fofbRecorder #(.BUFFER_CAPACITY(GPIO_RECORDER_CAPACITY),
               .CHANNEL_COUNT(GPIO_CHANNEL_COUNT),
               .DEBUG("false"))
  fofbRecorder (
    .clk(sysClk),
    .GPIO_OUT(GPIO_OUT),
    .csrStrobe(GPIO_STROBES[GPIO_IDX_WFR_CSR]),
    .pretriggerInitStrobe(GPIO_STROBES[GPIO_IDX_WFR_W_PRETRIGGER]),
    .posttriggerInitStrobe(GPIO_STROBES[GPIO_IDX_WFR_W_POSTTRIGGER]),
    .channelMapStrobe(GPIO_STROBES[GPIO_IDX_WFR_W_CHANNEL_BITMAP]),
    .addressStrobe(GPIO_STROBES[GPIO_IDX_WFR_ADDRESS]),
    .timestamp(sysTimestamp),
    .status(GPIO_IN[GPIO_IDX_WFR_CSR]),
    .triggerAddress(GPIO_IN[GPIO_IDX_WFR_ADDRESS]),
    .txData(GPIO_IN[GPIO_IDX_WFR_R_TX_DATA]),
    .rxData(GPIO_IN[GPIO_IDX_WFR_R_RX_DATA]),
    .acqTimestamp({GPIO_IN[GPIO_IDX_WFR_R_SECONDS],
                   GPIO_IN[GPIO_IDX_WFR_R_TICKS]}),
    .evrTrigger(evrTriggerBus[3]),
    .awgRunning(GPIO_IN[GPIO_IDX_AWG_CSR][29]),
    .tx_S_AXIS_TVALID(PS_SETPOINT_AXIS_TVALID),
    .tx_S_AXIS_TDATA(PS_SETPOINT_AXIS_TDATA),
    .tx_S_AXIS_TLAST(PS_SETPOINT_AXIS_TLAST),
    .rx_S_AXIS_TVALID(PS_READBACK_AXIS_TVALID),
    .rx_S_AXIS_TDATA(PS_READBACK_AXIS_TDATA),
    .rx_S_AXIS_TUSER(PS_READBACK_AXIS_TUSER));

//////////////////////////////////////////////////////////////////////////////
// Errant Electron Beam Interlock
eebi #(.SYSCLK_RATE(SYSCLK_RATE), .dbg("false")) eebi (
            .sysClk(sysClk),
            .sysCsrStrobe(GPIO_STROBES[GPIO_IDX_EEBI_CSR]),
            .sysCsrWriteData(GPIO_OUT),
            .sysCsr(GPIO_IN[GPIO_IDX_EEBI_CSR]),
            .sysTimestamp(sysTimestamp),
            .sysMostRecentFaultTime({GPIO_IN[GPIO_IDX_EEBI_FAULT_TIME_SECONDS],
                                     GPIO_IN[GPIO_IDX_EEBI_FAULT_TIME_TICKS]}),
            .auroraUserClk(auroraUserClk),
            .auroraFAstrobe(auroraFAstrobe),
            .localBPMvalues(localBPMvalues),
            .localBPMvaluesVALID(localBPMvaluesVALID),
            .eebiRelay(INTLK_RELAY_CTL),
            .eebiResetButton_n(INTLK_RESET_BUTTON_N));

//////////////////////////////////////////////////////////////////////////////
// Convert value from integer nm to double precision mm
errorConvert errorConvert (
          .clk(sysClk),
          .writeStrobe(GPIO_STROBES[GPIO_IDX_ERROR_CONVERT_WDATA]),
          .writeData(GPIO_OUT),
          .csrStrobe(GPIO_STROBES[GPIO_IDX_ERROR_CONVERT_CSR]),
          .status(GPIO_IN[GPIO_IDX_ERROR_CONVERT_CSR]),
          .resultHi(GPIO_IN[GPIO_IDX_ERROR_CONVERT_RDATA_HI]),
          .resultLo(GPIO_IN[GPIO_IDX_ERROR_CONVERT_RDATA_LO]));

/////////////////////////////////////////////////////////////////////////////
// Frequency counters
localparam FREQ_COUNTERS_NUM = 7;
localparam FREQ_SEL_WIDTH = $clog2(FREQ_COUNTERS_NUM+1);
reg  [FREQ_SEL_WIDTH-1:0] frequencyMonitorSelect;
wire [29:0] measuredFrequency;
always @(posedge sysClk) begin
    if (GPIO_STROBES[GPIO_IDX_FREQUENCY_MONITOR_CSR])
        frequencyMonitorSelect <= GPIO_OUT[FREQ_SEL_WIDTH-1:0];
end
assign GPIO_IN[GPIO_IDX_FREQUENCY_MONITOR_CSR] = { 2'b0, measuredFrequency };
wire auRefClk;  // TODO FIXME
freq_multi_count #(
        .NF(FREQ_COUNTERS_NUM),  // number of frequency counters in a block
        .NG(1),  // number of frequency counter blocks
        .gw(4),  // Gray counter width
        .cw(1),  // macro-cycle counter width
        .rw($clog2(SYSCLK_RATE*4/3)), // reference counter width
        .uw(30)) // unknown counter width
  frequencyCounters(
    .unk_clk({
        ethernetRxClk, ethernetTxClk,
        auRefClk,
        ethRefClk125Buff,
        auroraUserClk, evrClk, sysClk}),
    .refclk(sysClk),
    .refMarker(evrTriggerBus[1]),  // 1 PPS marker from event system
    .addr(frequencyMonitorSelect),
    .frequency(measuredFrequency));

/////////////////////////////////////////////////////////////////////////////
// Front panel
assign FP_LED0_GRN = evrTriggerBus[0];
assign FP_LED0_RED = 1'b0;
wire   FP_LED1_STATE_RED, FP_LED1_STATE_YELLOW, FP_LED1_STATE_GREEN;
assign FP_LED1_STATE_RED = !CELL_CCW_AuroraCoreStatus_channel_up
                        && !CELL_CW_AuroraCoreStatus_channel_up;
assign FP_LED1_STATE_GREEN = CELL_CCW_AuroraCoreStatus_channel_up
                          && CELL_CW_AuroraCoreStatus_channel_up;
assign FP_LED1_STATE_YELLOW = !FP_LED1_STATE_RED && !FP_LED1_STATE_GREEN;
assign FP_LED1_GRN = FP_LED1_STATE_YELLOW || FP_LED1_STATE_GREEN;
assign FP_LED1_RED = FP_LED1_STATE_YELLOW || FP_LED1_STATE_RED;

wire   FP_LED2_STATE_RED, FP_LED2_STATE_YELLOW, FP_LED2_STATE_GREEN;
assign FP_LED2_STATE_RED = !BPM_CCW_AuroraCoreStatus_channel_up
                        && !BPM_CW_AuroraCoreStatus_channel_up;
assign FP_LED2_STATE_GREEN = BPM_CCW_AuroraCoreStatus_channel_up
                          && BPM_CW_AuroraCoreStatus_channel_up;
assign FP_LED2_STATE_YELLOW = !FP_LED2_STATE_RED && !FP_LED2_STATE_GREEN;
assign FP_LED2_GRN = FP_LED2_STATE_YELLOW || FP_LED2_STATE_GREEN;
assign FP_LED2_RED = FP_LED2_STATE_YELLOW || FP_LED2_STATE_RED;

/////////////////////////////////////////////////////////////////////////////
// Marble LEDs
assign MARBLE_LD16 = evrTriggerBus[0];
assign MARBLE_LD17 = qsfp_led;

/////////////////////////////////////////////////////////////////////////////
// Miscellaneous
//`include "firmwareBuildDate.v"
assign GPIO_IN[GPIO_IDX_FIRMWARE_BUILD_DATE] = 0; // Deprecating firmware build date
`include "gitHash.vh"
assign GPIO_IN[GPIO_IDX_GITHASH] = GIT_REV_32BIT; // Deprecating firmware build date

/////////////////////////////////////////////////////////////////////////////
// FIFO/UART console I/O
fifoUART #(.CLK_RATE(SYSCLK_RATE),
           .BIT_RATE(115200)) fifoUART (
                   .clk(sysClk),
                   .strobe(GPIO_STROBES[GPIO_IDX_UART_CSR]),
                   .control(GPIO_OUT),
                   .status(GPIO_IN[GPIO_IDX_UART_CSR]),
                   .TxData(FPGA_RxD),
                   .RxData(FPGA_TxD));

//////////////////////////////////////////////////////////////////////////////
// Badger Ethernet MAC Interface
badger badger_i (
  .sysClk         (sysClk),  // TODO correct?
  .sysGPIO_OUT    (GPIO_OUT), // [31:0]
  .sysConfigStrobe(GPIO_STROBES[GPIO_IDX_NET_CONFIG_CSR]),
  .sysTxStrobe    (GPIO_STROBES[GPIO_IDX_NET_TX_CSR]),
  .sysRxStrobe    (GPIO_STROBES[GPIO_IDX_NET_RX_CSR]),
  .sysRxDataStrobe(GPIO_STROBES[GPIO_IDX_NET_RX_DATA]),
  .sysTxStatus    (GPIO_IN[GPIO_IDX_NET_TX_CSR]), // [31:0]
  .sysRxStatus    (GPIO_IN[GPIO_IDX_NET_RX_CSR]), // [31:0]
  .sysRxData      (GPIO_IN[GPIO_IDX_NET_RX_DATA]), // [31:0]

  // Two phases of 125 MHz clock, created by on-board reference
  .refClk125      (badgerRefClk125),
  .refClk125d90   (badgerRefClk125d90),

  // Diagnostic outputs (e.g. to frequency counters)
  .rx_clk(ethernetRxClk),
  .tx_clk(ethernetTxClk),

  // RGMII pins
  .RGMII_RX_CLK   (RGMII_RX_CLK),
  .RGMII_RX_CTRL  (RGMII_RX_CTRL),
  .RGMII_RXD      (RGMII_RXD), // [3:0]
  .RGMII_TX_CLK   (RGMII_TX_CLK),
  .RGMII_TX_CTRL  (RGMII_TX_CTRL),
  .RGMII_TXD      (RGMII_TXD) // [3:0]
);

`ifndef SIMULATE

//////////////////////////////////////////////////////////////////////////////
// Block design (MicroBlaze)

wire DUMMY_UART_LOOPBACK;

  system_marble system_i (
        .clkIn125(clkIn125), // input
        .badgerClk125(badgerRefClk125), // output
        .badgerClk125d90(badgerRefClk125d90), // output
        .clk200(clk200),  // output
        .sysClk(sysClk), // output
        .sysReset_n(sysReset_n),

        .auroraUserClk(auroraUserClk),
        .gt0_qplllock_out(gt0_qplllock_out),
        .gt0_qpllrefclklost_out(gt0_qpllrefclklost_out),
        .pll_not_locked_out(pll_not_locked_out),
        .auroraReset(auroraReset),
        .auroraRefClk(auRefClk),
        .gtxReset(sysGTXreset),
        .gtxResetOut(gtxResetOut),

        //.GT_DIFF_REFCLK_312_3_clk_n(MGT_CLK_1_N),
        //.GT_DIFF_REFCLK_312_3_clk_p(MGT_CLK_1_P),
        .GT_DIFF_REFCLK_125_clk_n(MGT_CLK_1_N),
        .GT_DIFF_REFCLK_125_clk_p(MGT_CLK_1_P),

        .BPM_CCW_AXI_STREAM_RX_tdata(BPM_CCW_AXI_STREAM_RX_tdata),
        .BPM_CCW_AXI_STREAM_RX_tlast(BPM_CCW_AXI_STREAM_RX_tlast),
        .BPM_CCW_AXI_STREAM_RX_tvalid(BPM_CCW_AXI_STREAM_RX_tvalid),
        .BPM_CCW_AuroraCoreStatus_channel_up(BPM_CCW_AuroraCoreStatus_channel_up),
        .BPM_CCW_AuroraCoreStatus_crc_pass_fail(BPM_CCW_AuroraCoreStatus_crc_pass_fail),
        .BPM_CCW_AuroraCoreStatus_crc_valid(BPM_CCW_AuroraCoreStatus_crc_valid),
        .BPM_CCW_AuroraCoreStatus_frame_err(BPM_CCW_AuroraCoreStatus_frame_err),
        .BPM_CCW_AuroraCoreStatus_hard_err(BPM_CCW_AuroraCoreStatus_hard_err),
        .BPM_CCW_AuroraCoreStatus_lane_up(BPM_CCW_AuroraCoreStatus_lane_up),
        .BPM_CCW_AuroraCoreStatus_rx_resetdone_out(BPM_CCW_AuroraCoreStatus_rx_resetdone_out),
        .BPM_CCW_AuroraCoreStatus_soft_err(BPM_CCW_AuroraCoreStatus_soft_err),
        .BPM_CCW_AuroraCoreStatus_tx_lock(BPM_CCW_AuroraCoreStatus_tx_lock),
        .BPM_CCW_AuroraCoreStatus_tx_resetdone_out(BPM_CCW_AuroraCoreStatus_tx_resetdone_out),
        .BPM_CCW_GT_RX_rxn(QSFP1_RX_N[1]),
        .BPM_CCW_GT_RX_rxp(QSFP1_RX_P[1]),
        .BPM_CCW_GT_TX_txn(QSFP1_TX_N[1]),
        .BPM_CCW_GT_TX_txp(QSFP1_TX_P[1]),

        .BPM_CW_AXI_STREAM_RX_tdata(BPM_CW_AXI_STREAM_RX_tdata),
        .BPM_CW_AXI_STREAM_RX_tlast(BPM_CW_AXI_STREAM_RX_tlast),
        .BPM_CW_AXI_STREAM_RX_tvalid(BPM_CW_AXI_STREAM_RX_tvalid),
        .BPM_CW_AuroraCoreStatus_channel_up(BPM_CW_AuroraCoreStatus_channel_up),
        .BPM_CW_AuroraCoreStatus_crc_pass_fail(BPM_CW_AuroraCoreStatus_crc_pass_fail),
        .BPM_CW_AuroraCoreStatus_crc_valid(BPM_CW_AuroraCoreStatus_crc_valid),
        .BPM_CW_AuroraCoreStatus_frame_err(BPM_CW_AuroraCoreStatus_frame_err),
        .BPM_CW_AuroraCoreStatus_hard_err(BPM_CW_AuroraCoreStatus_hard_err),
        .BPM_CW_AuroraCoreStatus_lane_up(BPM_CW_AuroraCoreStatus_lane_up),
        .BPM_CW_AuroraCoreStatus_rx_resetdone_out(BPM_CW_AuroraCoreStatus_rx_resetdone_out),
        .BPM_CW_AuroraCoreStatus_soft_err(BPM_CW_AuroraCoreStatus_soft_err),
        .BPM_CW_AuroraCoreStatus_tx_lock(BPM_CW_AuroraCoreStatus_tx_lock),
        .BPM_CW_AuroraCoreStatus_tx_resetdone_out(BPM_CW_AuroraCoreStatus_tx_resetdone_out),
        .BPM_CW_GT_RX_rxn(QSFP1_RX_N[2]),
        .BPM_CW_GT_RX_rxp(QSFP1_RX_P[2]),
        .BPM_CW_GT_TX_txn(QSFP1_TX_N[2]),
        .BPM_CW_GT_TX_txp(QSFP1_TX_P[2]),

        .CELL_CCW_AXI_STREAM_TX_tdata(CELL_CCW_AXI_STREAM_TX_tdata),
        .CELL_CCW_AXI_STREAM_TX_tlast(CELL_CCW_AXI_STREAM_TX_tlast),
        .CELL_CCW_AXI_STREAM_TX_tvalid(CELL_CCW_AXI_STREAM_TX_tvalid),
        .CELL_CCW_AXI_STREAM_TX_tready(CELL_CCW_AXI_STREAM_TX_tready),
        .CELL_CCW_AXI_STREAM_RX_tdata(CELL_CCW_AXI_STREAM_RX_tdata),
        .CELL_CCW_AXI_STREAM_RX_tlast(CELL_CCW_AXI_STREAM_RX_tlast),
        .CELL_CCW_AXI_STREAM_RX_tvalid(CELL_CCW_AXI_STREAM_RX_tvalid),
        .CELL_CCW_AuroraCoreStatus_channel_up(CELL_CCW_AuroraCoreStatus_channel_up),
        .CELL_CCW_AuroraCoreStatus_crc_pass_fail(CELL_CCW_AuroraCoreStatus_crc_pass_fail),
        .CELL_CCW_AuroraCoreStatus_crc_valid(CELL_CCW_AuroraCoreStatus_crc_valid),
        .CELL_CCW_AuroraCoreStatus_frame_err(CELL_CCW_AuroraCoreStatus_frame_err),
        .CELL_CCW_AuroraCoreStatus_hard_err(CELL_CCW_AuroraCoreStatus_hard_err),
        .CELL_CCW_AuroraCoreStatus_lane_up(CELL_CCW_AuroraCoreStatus_lane_up),
        .CELL_CCW_AuroraCoreStatus_rx_resetdone_out(CELL_CCW_AuroraCoreStatus_rx_resetdone_out),
        .CELL_CCW_AuroraCoreStatus_soft_err(CELL_CCW_AuroraCoreStatus_soft_err),
        .CELL_CCW_AuroraCoreStatus_tx_lock(CELL_CCW_AuroraCoreStatus_tx_lock),
        .CELL_CCW_AuroraCoreStatus_tx_resetdone_out(CELL_CCW_AuroraCoreStatus_tx_resetdone_out),
        .CELL_CCW_GT_RX_rxn(QSFP2_RX_N[0]),
        .CELL_CCW_GT_RX_rxp(QSFP2_RX_P[0]),
        .CELL_CCW_GT_TX_txn(QSFP2_TX_N[0]),
        .CELL_CCW_GT_TX_txp(QSFP2_TX_P[0]),

        .CELL_CW_AXI_STREAM_TX_tdata(CELL_CW_AXI_STREAM_TX_tdata),
        .CELL_CW_AXI_STREAM_TX_tlast(CELL_CW_AXI_STREAM_TX_tlast),
        .CELL_CW_AXI_STREAM_TX_tvalid(CELL_CW_AXI_STREAM_TX_tvalid),
        .CELL_CW_AXI_STREAM_TX_tready(CELL_CW_AXI_STREAM_TX_tready),
        .CELL_CW_AXI_STREAM_RX_tdata(CELL_CW_AXI_STREAM_RX_tdata),
        .CELL_CW_AXI_STREAM_RX_tlast(CELL_CW_AXI_STREAM_RX_tlast),
        .CELL_CW_AXI_STREAM_RX_tvalid(CELL_CW_AXI_STREAM_RX_tvalid),
        .CELL_CW_AuroraCoreStatus_channel_up(CELL_CW_AuroraCoreStatus_channel_up),
        .CELL_CW_AuroraCoreStatus_crc_pass_fail(CELL_CW_AuroraCoreStatus_crc_pass_fail),
        .CELL_CW_AuroraCoreStatus_crc_valid(CELL_CW_AuroraCoreStatus_crc_valid),
        .CELL_CW_AuroraCoreStatus_frame_err(CELL_CW_AuroraCoreStatus_frame_err),
        .CELL_CW_AuroraCoreStatus_hard_err(CELL_CW_AuroraCoreStatus_hard_err),
        .CELL_CW_AuroraCoreStatus_lane_up(CELL_CW_AuroraCoreStatus_lane_up),
        .CELL_CW_AuroraCoreStatus_rx_resetdone_out(CELL_CW_AuroraCoreStatus_rx_resetdone_out),
        .CELL_CW_AuroraCoreStatus_soft_err(CELL_CW_AuroraCoreStatus_soft_err),
        .CELL_CW_AuroraCoreStatus_tx_lock(CELL_CW_AuroraCoreStatus_tx_lock),
        .CELL_CW_AuroraCoreStatus_tx_resetdone_out(CELL_CW_AuroraCoreStatus_tx_resetdone_out),
        .CELL_CW_GT_RX_rxn(QSFP2_RX_N[1]),
        .CELL_CW_GT_RX_rxp(QSFP2_RX_P[1]),
        .CELL_CW_GT_TX_txn(QSFP2_TX_N[1]),
        .CELL_CW_GT_TX_txp(QSFP2_TX_P[1]),

        .evr_mgt_rec_clk(evrClk),
        .evr_mgt_par_data(evr_mgt_par_data & {16{evrRxLocked}}),
        .evr_mgt_chariscomma(evr_mgt_chariscomma),
        .evr_mgt_charisk(evr_mgt_charisk),
        .evr_mgt_reset_done(evr_mgt_reset_done),
        .evrTriggerBus(evrTriggerBus),
        .evrDataBus(evrDataBus),
        .evrTimestamp(evrTimestamp),
        .evr_mgt_drp_daddr(evr_mgt_drp_daddr),
        .evr_mgt_drp_den(evr_mgt_drp_den),
        .evr_mgt_drp_di(evr_mgt_drp_di),
        .evr_mgt_drp_do(evr_mgt_drp_do),
        .evr_mgt_drp_drdy(evr_mgt_drp_drdy),
        .evr_mgt_drp_dwe(evr_mgt_drp_dwe),

        .BRAM_BPM_SETPOINTS_ADDR(BRAM_BPM_SETPOINTS_ADDR),
        .BRAM_BPM_SETPOINTS_WDATA(BRAM_BPM_SETPOINTS_WDATA),
        .BRAM_BPM_SETPOINTS_WENABLE(BRAM_BPM_SETPOINTS_WENABLE),
        .BRAM_BPM_SETPOINTS_RDATA(BRAM_BPM_SETPOINTS_RDATA),

        // Dummy UART to keep SDK tools happy
        .uart_rtl_rxd(DUMMY_UART_LOOPBACK),
        .uart_rtl_txd(DUMMY_UART_LOOPBACK),

        .GPIO_IN(GPIO_IN_FLATTENED),
        .GPIO_OUT(GPIO_OUT),
        .GPIO_STROBES(GPIO_STROBES));
`endif // `ifndef SIMULATE

endmodule
