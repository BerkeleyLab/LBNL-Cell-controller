localparam GIT_REV_STR = "8824da04";
localparam GIT_DIRTY = 1;
localparam GIT_REV_32BIT = 32'h8824da04;
